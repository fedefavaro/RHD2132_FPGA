-----------------------------------------------------------------------------------------------------------------------
-- Author:
-- 
-- Create Date:		13/11/2016  -- dd/mm/yyyy
-- Module Name:		test_maquina_control
-- Project Name:
-- Target Devices:
-- Tool versions:
-- Description: 
--
--		...
--      
-----------------------------------------------------------------------------------------------------------------------

LIBRARY ieee ;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;


ENTITY test_maquina_control IS
       PORT(
          CLK                       : IN  STD_LOGIC;
          RESET                     : IN  STD_LOGIC;
          -- registros param chips --
          
          -- registros control --
          
       );
END test_maquina_control;


ARCHITECTURE synth of test_maquina_control IS


BEGIN



END synth;


